

module our;
	initial begin
		$display("hello again, world");
		$finish;
	end
endmodule





















